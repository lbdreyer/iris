dimensions:
	dim0 = 10 ;
variables:
	double temp(dim0) ;
		temp:standard_name = "air_temperature" ;
		temp:units = "K" ;
		temp:coordinates = "time" ;
	int64 time(dim0) ;
		time:units = "1" ;
		time:standard_name = "time" ;
	double temp3(dim0) ;
		temp3:long_name = "air_temperature" ;
		temp3:units = "K" ;
		temp3:coordinates = "time_0" ;
	int64 time_0(dim0) ;
		time_0:units = "1" ;
		time_0:standard_name = "time" ;

// global attributes:
		:Conventions" = "CF-1.7" ;
}
